`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 21.04.2023 23:53:47
// Design Name: 
// Module Name: simulation
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module simulation(
    
    );
//    reg clk;
//    reg grant_line;
//    wire [12:0] hit_counter;
//    wire [20:0] counter;
//    initial 
//    begin
//        grant_line=0;
//        clk=1;
//        forever
//        #1 clk=~clk;
//    end
//    reg [31:0] address;
    
//    wire [31:0] done_address;
//    wire done;
////    wire [19:0] out_counter;
//    Memory mem(.clk(clk),.address(address),.grant_line(grant_line),.done_address(done_address),.done(done),.hit_counter(hit_counter),.counter(counter));
//    initial
//    begin
//        grant_line=1; address= 10;
//        #2 grant_line=0;
//        #18 grant_line=1; address= 2048;
//        #2 grant_line=0;
//        #18 grant_line=1; address= 2049;
//        #2 grant_line=0;
//        #18 grant_line=1; address= 2050;
//        #2 grant_line=0;
//        #18 grant_line=1; address= 10;
//        #2 grant_line=0;
////        #18 grant_line=1; address= 10;
////        #2 grant_line=0;
////        #18 grant_line=1; address= 10;
////        #2 grant_line=0;
////        #18 grant_line=1; address= 10;
////        #2 grant_line=0;
////        #18 grant_line=1; address= 10;
////        #2 grant_line=0;
////        #18 grant_line=1; address= 10;
////        #2 grant_line=0;
////        #18 grant_line=1; address= 10;
////        #2 grant_line=0;
////        #18 grant_line=1; address= 10;
////        #2 grant_line=0;
        
//        #400;
//    end
reg clk;
//reg en;
//reg iamtaking;
reg [31:0] data_in;
reg en;
//reg [31:0] mem_ins;
//reg recieved;
//wire [31:0] data_out;
//wire iamsending;
wire[12:0] hit_counter;
wire[12:0] miss_counter;
wire[20:0] counter;


initial
    begin
//        en=0;
        clk=1;
        en=0;
//        iamtaking=0;
//        recieved=0;
        forever
        #1 clk=~clk;
    end

top t(clk,data_in,en,hit_counter,counter);

initial 
begin
//data_in=1;
//#2 data_in=2;
//#2 data_in=3;
//#2 data_in=2;
//#2 data_in=4;
//#2 data_in=2048;
//#2 data_in=5;
//#2 data_in=6;
//#2 data_in=2049;
//#2 data_in=19;
//#2 data_in=20;
//#2 data_in=21;

 data_in='h00004138 ;
#2 data_in='h00004140 ;
#2 data_in='h00002866 ;
#2 data_in='h00002882 ;
#2 data_in='h00005664 ;
#2 data_in='h00002cc1 ;
#2 data_in='h0000297e ;
#2 data_in='h00002982 ;
#2 data_in='h00003535 ;
#2 data_in='h00006214 ;
#2 data_in='h0000446b ;
#2 data_in='h00004483 ;
#2 data_in='h00004d65 ;
#2 data_in='h000033dc ;
#2 data_in='h0000739d ;
#2 data_in='h000047ec ;
#2 data_in='h000026ea ;
#2 data_in='h000058af ;
#2 data_in='h000058c3 ;
#2 data_in='h00005e06 ;
#2 data_in='h00004873 ;
#2 data_in='h00004643 ;
#2 data_in='h00006ce4 ;
#2 data_in='h00006d00 ;
#2 data_in='h00004e06 ;
#2 data_in='h000037e4 ;
#2 data_in='h00003e85 ;
#2 data_in='h0000375c ;
#2 data_in='h00003780 ;
#2 data_in='h00007b8d ;
#2 data_in='h0000427b ;
#2 data_in='h00004283 ;
#2 data_in='h0000545f ;
#2 data_in='h00005364 ;
#2 data_in='h0000773f ;
#2 data_in='h0000551a ;
#2 data_in='h0000616e ;
#2 data_in='h00004b0e ;
#2 data_in='h000036cd ;
#2 data_in='h000029c1 ;
#2 data_in='h00006bce ;
#2 data_in='h000070ef ;
#2 data_in='h00007103 ;
#2 data_in='h00002542 ;
#2 data_in='h00004920 ;
#2 data_in='h000079e9 ;
#2 data_in='h000065e4 ;
#2 data_in='h00006da4 ;
#2 data_in='h00007dc3 ;
#2 data_in='h0000478e ;
#2 data_in='h000072c1 ;
#2 data_in='h00003430 ;
#2 data_in='h00002d7c ;
#2 data_in='h00002d80 ;
#2 data_in='h000062bb ;
#2 data_in='h00007763 ;
#2 data_in='h0000332d ;
#2 data_in='h00007ea2 ;
#2 data_in='h000022b1 ;
#2 data_in='h00006280 ;
#2 data_in='h00005a55 ;
#2 data_in='h00005037 ;
#2 data_in='h00006468 ;
#2 data_in='h00006480 ;
#2 data_in='h000054ea ;
#2 data_in='h00004b85 ;
#2 data_in='h00002fdd ;
#2 data_in='h000022ef ;
#2 data_in='h00004e4e ;
#2 data_in='h000070a2 ;
#2 data_in='h000043a7 ;
#2 data_in='h0000706b ;
#2 data_in='h00005b2b ;
#2 data_in='h00007626 ;
#2 data_in='h0000577a ;
#2 data_in='h00004545 ;
#2 data_in='h00006874 ;
#2 data_in='h000061ff ;
#2 data_in='h00003ac7 ;
#2 data_in='h000076c6 ;
#2 data_in='h00005ef2 ;
#2 data_in='h000071fe ;
#2 data_in='h00004d2c ;
#2 data_in='h00005dff ;
#2 data_in='h00004730 ;
#2 data_in='h00004983 ;
#2 data_in='h00006c5f ;
#2 data_in='h000056cd ;
#2 data_in='h00007ac4 ;
#2 data_in='h00007c28 ;
#2 data_in='h00004426 ;
#2 data_in='h00004b42 ;
#2 data_in='h00003d96 ;
#2 data_in='h000035dc ;
#2 data_in='h000044f5 ;
#2 data_in='h0000698f ;
#2 data_in='h00003656 ;
#2 data_in='h00007e3f ;
#2 data_in='h00002b83 ;
#2 data_in='h00004f01 ;
#2 data_in='h000036ae ;
#2 data_in='h00006c83 ;
#2 data_in='h00003081 ;
#2 data_in='h0000798a ;
#2 data_in='h00003a99 ;
#2 data_in='h0000315b ;
#2 data_in='h00004af7 ;
#2 data_in='h000045d1 ;
#2 data_in='h000024e1 ;
#2 data_in='h00007d4e ;
#2 data_in='h0000790a ;
#2 data_in='h00006d70 ;
#2 data_in='h00003f52 ;
#2 data_in='h00007b75 ;
#2 data_in='h00003b91 ;
#2 data_in='h00003f99 ;
#2 data_in='h00005607 ;
#2 data_in='h000055a8 ;
#2 data_in='h00007425 ;
#2 data_in='h00005fb2 ;
#2 data_in='h00005ccc ;
#2 data_in='h00003042 ;
#2 data_in='h00002a49 ;
#2 data_in='h00002b08 ;
#2 data_in='h000046d2 ;
#2 data_in='h00003cc6 ;
#2 data_in='h00004f97 ;
#2 data_in='h00006517 ;
#2 data_in='h00005998 ;
#2 data_in='h00007a00 ;
#2 data_in='h00007c9e ;
#2 data_in='h00007cc2 ;
#2 data_in='h00006661 ;
#2 data_in='h00003196 ;
#2 data_in='h00007677 ;
#2 data_in='h0000640e ;
#2 data_in='h00007285 ;
#2 data_in='h0000394d ;
#2 data_in='h00005a2d ;
#2 data_in='h00002a01 ;
#2 data_in='h0000261e ;
#2 data_in='h000026d8 ;
#2 data_in='h00002700 ;
#2 data_in='h000067c0 ;
#2 data_in='h00004947 ;
#2 data_in='h00004fc2 ;
#2 data_in='h0000637d ;
#2 data_in='h00006381 ;
#2 data_in='h00004380 ;
#2 data_in='h000042ea ;
#2 data_in='h00004833 ;
#2 data_in='h00004aaf ;
#2 data_in='h000071a7 ;
#2 data_in='h00002c08 ;
#2 data_in='h00005d55 ;
#2 data_in='h000060d1 ;
#2 data_in='h00007825 ;
#2 data_in='h00005e8a ;
#2 data_in='h00005543 ;
#2 data_in='h00003c1b ;
#2 data_in='h00002c40 ;
#2 data_in='h000048a1 ;
#2 data_in='h00004625 ;
#2 data_in='h00003849 ;
#2 data_in='h00003d4b ;
#2 data_in='h00005d82 ;
#2 data_in='h00004efb ;
#2 data_in='h000021c7 ;
#2 data_in='h000061c0 ;
#2 data_in='h00005799 ;
#2 data_in='h000057c1 ;
#2 data_in='h00003e6f ;
#2 data_in='h00003b02 ;
#2 data_in='h00007ab5 ;
#2 data_in='h000069fb ;
#2 data_in='h00006a03 ;
#2 data_in='h00003d3a ;
#2 data_in='h00005bb5 ;
#2 data_in='h00005bc1 ;
#2 data_in='h00005fe7 ;
#2 data_in='h00003b42 ;
#2 data_in='h000051ff ;
#2 data_in='h00003dff ;
#2 data_in='h00003e03 ;
#2 data_in='h00004519 ;
#2 data_in='h00007245 ;
#2 data_in='h00007da1 ;
#2 data_in='h00006069 ;
#2 data_in='h00006081 ;
#2 data_in='h000054bf ;
#2 data_in='h00002dea ;
#2 data_in='h00006e36 ;
#2 data_in='h00002e14 ;
#2 data_in='h0000670c ;
#2 data_in='h000047e4 ;
#2 data_in='h00003ed6 ;
#2 data_in='h00003f02 ;
#2 data_in='h000063c2 ;
#2 data_in='h00002432 ;
#2 data_in='h000046aa ;
#2 data_in='h00005957 ;
#2 data_in='h00006338 ;
#2 data_in='h00005278 ;
#2 data_in='h00007f6a ;
#2 data_in='h00006815 ;
#2 data_in='h0000402d ;
#2 data_in='h00004041 ;
#2 data_in='h00006b52 ;
#2 data_in='h000062b0 ;
#2 data_in='h00002280 ;
#2 data_in='h00007244 ;
#2 data_in='h00004ce2 ;
#2 data_in='h00005642 ;
#2 data_in='h00003831 ;
#2 data_in='h0000221e ;
#2 data_in='h00006881 ;
#2 data_in='h00007b1e ;
#2 data_in='h00004737 ;
#2 data_in='h00004743 ;
#2 data_in='h00002321 ;
#2 data_in='h00004c8d ;
#2 data_in='h00005386 ;
#2 data_in='h00003fde ;
#2 data_in='h00005e78 ;
#2 data_in='h00004230 ;
#2 data_in='h000052dc ;
#2 data_in='h00002241 ;
#2 data_in='h00006593 ;
#2 data_in='h00006961 ;
#2 data_in='h00002b70 ;
#2 data_in='h00007325 ;
#2 data_in='h0000542a ;
#2 data_in='h00006ea3 ;
#2 data_in='h00002ee3 ;
#2 data_in='h00005f22 ;
#2 data_in='h0000652c ;
#2 data_in='h000032fc ;
#2 data_in='h00007a59 ;
#2 data_in='h00006dc7 ;
#2 data_in='h00005d12 ;
#2 data_in='h00006260 ;
#2 data_in='h00002240 ;
#2 data_in='h00005703 ;
#2 data_in='h000075a6 ;
#2 data_in='h00002948 ;
#2 data_in='h00006ab4 ;
#2 data_in='h00004a53 ;
#2 data_in='h00005cb4 ;
#2 data_in='h00004ab5 ;
#2 data_in='h000040b6 ;
#2 data_in='h00006080 ;
#2 data_in='h000040c2 ;
#2 data_in='h000060c0 ;
#2 data_in='h00002725 ;
#2 data_in='h00007861 ;
#2 data_in='h00007881 ;
#2 data_in='h0000581d ;
#2 data_in='h00002bf9 ;
#2 data_in='h00002371 ;
#2 data_in='h0000398f ;
#2 data_in='h000039c3 ;
#2 data_in='h00005856 ;
#2 data_in='h00006110 ;
#2 data_in='h00004100 ;
#2 data_in='h00002078 ;
#2 data_in='h00006040 ;
#2 data_in='h00002080 ;
#2 data_in='h00004080 ;
#2 data_in='h000078fd ;
#2 data_in='h00002659 ;
#2 data_in='h00007972 ;
#2 data_in='h000020c4 ;
#2 data_in='h00007bd1 ;
#2 data_in='h000031c3 ;
#2 data_in='h000060c9 ;
#2 data_in='h000020c0 ;
#2 data_in='h00002683 ;
#2 data_in='h000053ea ;
#2 data_in='h00003c4c ;
#2 data_in='h00003bf4 ;
#2 data_in='h00004c4e ;
#2 data_in='h000028da ;
#2 data_in='h00003936 ;
#2 data_in='h00005b66 ;
#2 data_in='h0000591b ;
#2 data_in='h000033a3 ;
#2 data_in='h000027b0 ;
#2 data_in='h00003f3a ;
#2 data_in='h000071fe ;
#2 data_in='h00007202 ;
#2 data_in='h0000523c ;
#2 data_in='h00006f10 ;
#2 data_in='h00007bd9 ;
#2 data_in='h00004bc1 ;
#2 data_in='h00005068 ;
#2 data_in='h00005080 ;
#2 data_in='h0000690b ;
#2 data_in='h00003621 ;
#2 data_in='h00005a97 ;
#2 data_in='h000035bb ;
#2 data_in='h00002503 ;
#2 data_in='h00005fc2 ;
#2 data_in='h00006e41 ;
#2 data_in='h00006c01 ;
#2 data_in='h00003ca7 ;
#2 data_in='h0000246c ;
#2 data_in='h00002480 ;
#2 data_in='h00002cb3 ;
#2 data_in='h0000675f ;
#2 data_in='h000030dd ;
#2 data_in='h00004a16 ;
#2 data_in='h00002740 ;
#2 data_in='h0000716f ;
#2 data_in='h000023e7 ;
#2 data_in='h000051cb ;
#2 data_in='h000067ba ;
#2 data_in='h00002e9e ;
#2 data_in='h000051bf ;
#2 data_in='h00003480 ;
#2 data_in='h00007e6c ;
#2 data_in='h0000342f ;
#2 data_in='h00002aa5 ;
#2 data_in='h00002ac1 ;
#2 data_in='h00004334 ;
#2 data_in='h00004340 ;
#2 data_in='h00006340 ;
#2 data_in='h00007452 ;
#2 data_in='h00005c55 ;
#2 data_in='h00003525 ;
#2 data_in='h00005f2e ;
#2 data_in='h000066fd ;
#2 data_in='h000034c6 ;
#2 data_in='h00007778 ;
#2 data_in='h00007780 ;
#2 data_in='h000068c3 ;
#2 data_in='h000045b3 ;
#2 data_in='h00006012 ;
#2 data_in='h00004000 ;
#2 data_in='h0000320f ;
#2 data_in='h00003342 ;
#2 data_in='h00005ada ;
#2 data_in='h00006a6b ;
#2 data_in='h00007c68 ;
#2 data_in='h00007541 ;
#2 data_in='h00004e81 ;
#2 data_in='h00005202 ;
#2 data_in='h00003001 ;
#2 data_in='h00007d1a ;
#2 data_in='h0000737f ;
#2 data_in='h000076bf ;
#2 data_in='h00007703 ;
#2 data_in='h00007ec3 ;
#2 data_in='h00006f47 ;
#2 data_in='h000041a8 ;
#2 data_in='h00003fbb ;
#2 data_in='h0000213e ;
#2 data_in='h00006100 ;
#2 data_in='h00002142 ;
#2 data_in='h00006140 ;
#2 data_in='h00007483 ;
#2 data_in='h000062d0 ;
#2 data_in='h000022c0 ;
#2 data_in='h00002f6c ;
#2 data_in='h00006ee9 ;
#2 data_in='h000052a6 ;
#2 data_in='h0000696b ;
#2 data_in='h00005130 ;
#2 data_in='h00005432 ;
#2 data_in='h00005300 ;
#2 data_in='h00006775 ;
#2 data_in='h000066a3 ;
#2 data_in='h000049c0 ;
#2 data_in='h00005f66 ;
#2 data_in='h00007e29 ;
#2 data_in='h00002d03 ;
#2 data_in='h0000494c ;
#2 data_in='h00005169 ;
#2 data_in='h0000604e ;
#2 data_in='h00004040 ;
#2 data_in='h0000324d ;
#2 data_in='h000059f0 ;
#2 data_in='h000075f4 ;
#2 data_in='h000046db ;
#2 data_in='h0000370c ;
#2 data_in='h00003456 ;
#2 data_in='h000034bd ;
#2 data_in='h00007fec ;
#2 data_in='h00008000 ;
#2 data_in='h00002d7a ;
#2 data_in='h000048e6 ;
#2 data_in='h000027d0 ;
#2 data_in='h00003886 ;
#2 data_in='h000025e0 ;
#2 data_in='h00002037 ;
#2 data_in='h00006000 ;
#2 data_in='h00003355 ;
#2 data_in='h000032be ;
#2 data_in='h00003a39 ;
#2 data_in='h000064c1 ;
#2 data_in='h0000611d ;
#2 data_in='h00002100 ;
#2 data_in='h00002e45 ;
#2 data_in='h0000401c ;
#2 data_in='h00008000 ;
#2 data_in='h00004040 ;
#2 data_in='h00007f4b ;
#2 data_in='h00006fff ;
#2 data_in='h00004d93 ;
#2 data_in='h00003125 ;
#2 data_in='h00007f31 ;
#2 data_in='h00006b8c ;
#2 data_in='h000073fe ;
#2 data_in='h00003574 ;
#2 data_in='h000050de ;
#2 data_in='h00002583 ;
#2 data_in='h00006080 ;
#2 data_in='h000041d9 ;
#2 data_in='h000023ac ;
#2 data_in='h00002800 ;
#2 data_in='h000071fb ;
#2 data_in='h00003642 ;
#2 data_in='h000077f2 ;
#2 data_in='h000043d8 ;
#2 data_in='h00004083 ;
#2 data_in='h00002080 ;
#2 data_in='h0000603a ;
#2 data_in='h00004000 ;
#2 data_in='h00004381 ;
#2 data_in='h000022d4 ;
#2 data_in='h000042c0 ;
#2 data_in='h00006342 ;
#2 data_in='h00004340 ;
#2 data_in='h000020f1 ;
#2 data_in='h00002101 ;
#2 data_in='h00006518 ;
#2 data_in='h000033cb ;
#2 data_in='h0000410a ;
#2 data_in='h00006100 ;
#2 data_in='h00004c1c ;
#2 data_in='h00007000 ;
#2 data_in='h000042fb ;
#2 data_in='h000062c0 ;
#2 data_in='h000055da ;
#2 data_in='h0000617c ;
#2 data_in='h00004140 ;
#2 data_in='h00006180 ;
#2 data_in='h000062e2 ;
#2 data_in='h000022c0 ;
#2 data_in='h00002180 ;
#2 data_in='h00004de8 ;
#2 data_in='h00006b26 ;
#2 data_in='h00006105 ;
#2 data_in='h00002100 ;
#2 data_in=-1;
#2 en = 1;
$finish;
end

endmodule